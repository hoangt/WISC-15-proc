module pipeline_control();
//TODO: Determine what control signals are needed at each level to determine a stall.
endmodule
